package version_pkg;
  // Other declarations can go here...

  // Auto-updated version and date constants
  localparam logic [7:0]  C_VERSION_MAJOR  = 8'd0;
  localparam logic [7:0]  C_VERSION_MINOR  = 8'd0;
  localparam logic [7:0]  C_VERSION_PATCH  = 8'd0;
  localparam logic [7:0]  C_VERSION_BUILD  = 8'd77;

  localparam logic [15:0] C_VERSION_YEAR   = 16'h2026;
  localparam logic [7:0]  C_VERSION_MONTH  = 8'h01;
  localparam logic [7:0]  C_VERSION_DAY    = 8'h15;
  localparam logic [7:0]  C_VERSION_HOUR   = 8'h12;
  localparam logic [7:0]  C_VERSION_MINUTE = 8'h15;
  localparam logic [7:0]  C_VERSION_SECOND = 8'h48;

endpackage : version_pkg
