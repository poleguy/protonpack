package version_pkg;
  // Other declarations can go here...

  // Auto-updated version and date constants
  localparam logic [7:0]  C_VERSION_MAJOR  = 8'd0;
  localparam logic [7:0]  C_VERSION_MINOR  = 8'd0;
  localparam logic [7:0]  C_VERSION_PATCH  = 8'd0;
  localparam logic [7:0]  C_VERSION_BUILD  = 8'd53;

  localparam logic [15:0] C_VERSION_YEAR   = 16'h2025;
  localparam logic [7:0]  C_VERSION_MONTH  = 8'h11;
  localparam logic [7:0]  C_VERSION_DAY    = 8'h05;
  localparam logic [7:0]  C_VERSION_HOUR   = 8'h13;
  localparam logic [7:0]  C_VERSION_MINUTE = 8'h55;
  localparam logic [7:0]  C_VERSION_SECOND = 8'h09;

endpackage : version_pkg
