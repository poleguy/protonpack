obsolete, use verilog version.