------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gt_serial_telem_rx_subsystem.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module gt_serial_telem_rx_subsystem
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned."+";

library UNISIM;
use UNISIM.VCOMPONENTS.all;

library work;
use work.telemetry_cfg_pkg.all;

--library xil_defaultlib;
--use xil_defaultlib.all;

--***********************************Entity Declaration************************

entity gt_serial_telem_rx_subsystem is
  generic
    (
      EXAMPLE_CONFIG_INDEPENDENT_LANES : integer   := 1;
      EXAMPLE_LANE_WITH_START_CHAR     : integer   := 0;  -- specifies lane with unique start frame ch
      EXAMPLE_WORDS_IN_BRAM            : integer   := 512;  -- specifies amount of data in BRAM
      EXAMPLE_SIM_GTRESET_SPEEDUP      : string    := "FALSE";  -- simulation setting for GT SecureIP model
      STABLE_CLOCK_PERIOD              : integer   := 7;
      EXAMPLE_USE_CHIPSCOPE            : integer   := 1;  -- Set to 1 to use Chipscope to drive resets
      g_debug                          : std_logic := '0'
      );
  port
    (
      Q0_CLK1_GTREFCLK_PAD_N_IN : in  std_logic; -- 125MHz
      Q0_CLK1_GTREFCLK_PAD_P_IN : in  std_logic;
      DRP_CLK_IN                : in  std_logic;  -- would be the 128Mhz coming direct from si570 (AS)
      rst_128M                  : in std_logic;
      -- GTTX_RESET_IN                           : in   std_logic;
      -- GTRX_RESET_IN                           : in   std_logic;
      -- PLL0_RESET_IN                           : in   std_logic; 
      -- PLL1_RESET_IN                           : in   std_logic;
--      TRACK_DATA_OUT            : out std_logic;
      SOFT_RESET_OUT            : out std_logic;
      RXN_IN                    : in  std_logic;
      RXP_IN                    : in  std_logic;
      TXN_OUT                   : out std_logic;
      TXP_OUT                   : out std_logic;
      -- 128MHz data out from recovered clock does not need a valid
      DATA_OUT                  : out std_logic_vector(31 downto 0); 
      DATA_CLK_OUT                  : out std_logic; 
      DATA_IS_K_OUT             : out std_logic_vector(3 downto 0)
      );


end gt_serial_telem_rx_subsystem;

architecture RTL of gt_serial_telem_rx_subsystem is
  attribute DowngradeIPIdentifiedWarnings        : string;
  attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

  attribute CORE_GENERATION_INFO        : string;
  attribute CORE_GENERATION_INFO of RTL : architecture is "gt_serial_telem_rx,gtwizard_v3_6_9,{protocol_file=Start_from_scratch}";

--**************************Component Declarations*****************************
--    component gt_serial_telem_rx
--        port
--        (
--            SOFT_RESET_TX_IN                        : in   std_logic;
--            SOFT_RESET_RX_IN                        : in   std_logic;
--            DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
--            Q0_CLK1_GTREFCLK_PAD_N_IN               : in   std_logic;
--            Q0_CLK1_GTREFCLK_PAD_P_IN               : in   std_logic;
--
--            GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
--            GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
--            GT0_DATA_VALID_IN                       : in   std_logic;
--            GT0_TX_MMCM_LOCK_OUT                    : out  std_logic;
--            GT0_RX_MMCM_LOCK_OUT                    : out  std_logic;
--         
--            GT0_TXUSRCLK_OUT                        : out  std_logic;
--            GT0_TXUSRCLK2_OUT                       : out  std_logic;
--            GT0_RXUSRCLK_OUT                        : out  std_logic;
--            GT0_RXUSRCLK2_OUT                       : out  std_logic;
--
--            --_________________________________________________________________________
--            --GT0  (X0Y3)
--            --____________________________CHANNEL PORTS________________________________
--            ---------------------------- Channel - DRP Ports  --------------------------
--            gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
--            gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
--            gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
--            gt0_drpen_in                            : in   std_logic;
--            gt0_drprdy_out                          : out  std_logic;
--            gt0_drpwe_in                            : in   std_logic;
--            --------------------- RX Initialization and Reset Ports --------------------
--            gt0_eyescanreset_in                     : in   std_logic;
--            gt0_rxuserrdy_in                        : in   std_logic;
--            -------------------------- RX Margin Analysis Ports ------------------------
--            gt0_eyescandataerror_out                : out  std_logic;
--            gt0_eyescantrigger_in                   : in   std_logic;
--            ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--            gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
--            ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
--            gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
--            gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
--            gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
--            ------------------------ Receive Ports - RX AFE Ports ----------------------
--            gt0_gtprxn_in                           : in   std_logic;
--            gt0_gtprxp_in                           : in   std_logic;
--            -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
--            gt0_rxslide_in                          : in   std_logic;
--            ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
--            gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
--            -------------------- Receive Ports - RX Equailizer Ports -------------------
--            gt0_rxlpmhfhold_in                      : in   std_logic;
--            gt0_rxlpmlfhold_in                      : in   std_logic;
--            --------------- Receive Ports - RX Fabric Output Control Ports -------------
--            gt0_rxoutclkfabric_out                  : out  std_logic;
--            ------------- Receive Ports - RX Initialization and Reset Ports ------------
--            gt0_gtrxreset_in                        : in   std_logic;
--            gt0_rxlpmreset_in                       : in   std_logic;
--            -------------- Receive Ports -RX Initialization and Reset Ports ------------
--            gt0_rxresetdone_out                     : out  std_logic;
--            --------------------- TX Initialization and Reset Ports --------------------
--            gt0_gttxreset_in                        : in   std_logic;
--            gt0_txuserrdy_in                        : in   std_logic;
--            ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--            gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
--            ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
--            gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);
--            --------------- Transmit Ports - TX Configurable Driver Ports --------------
--            gt0_gtptxn_out                          : out  std_logic;
--            gt0_gtptxp_out                          : out  std_logic;
--            ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--            gt0_txoutclkfabric_out                  : out  std_logic;
--            gt0_txoutclkpcs_out                     : out  std_logic;
--            ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--            gt0_txresetdone_out                     : out  std_logic;
--
--            --____________________________COMMON PORTS________________________________
--           GT0_PLL0RESET_OUT  : out std_logic;
--                 GT0_PLL0OUTCLK_OUT  : out std_logic;
--                          GT0_PLL0OUTREFCLK_OUT  : out std_logic;
--                                   GT0_PLL0LOCK_OUT  : out std_logic;
--                                            GT0_PLL0REFCLKLOST_OUT  : out std_logic;    
--                                                     GT0_PLL1OUTCLK_OUT  : out std_logic;
--                                                              GT0_PLL1OUTREFCLK_OUT  : out std_logic;
--
--                                                                      sysclk_in : in std_logic
--                                                                  );
--    end component;
--
--
--
--    component gt_serial_telem_rx_GT_FRAME_GEN 
--        generic
--        (
--             WORDS_IN_BRAM    : integer := 512
--         );
--        port
--        (
--            -- User Interface
--        TX_DATA_OUT             : out   std_logic_vector(79 downto 0);
--        TXCTRL_OUT              : out   std_logic_vector(7 downto 0); 
--            -- System Interface
--        USER_CLK                : in    std_logic;      
--        SYSTEM_RESET            : in    std_logic
--    ); 
--    end component;
--
--    component gt_serial_telem_rx_GT_FRAME_CHECK 
--        generic
--        (
--            RX_DATA_WIDTH            : integer := 16;
--            RXCTRL_WIDTH             : integer := 2; 
--            WORDS_IN_BRAM            : integer := 256;
--            CHANBOND_SEQ_LEN         : integer := 1;
--            COMMA_DOUBLE             : std_logic_vector(15 downto 0) := x"f628";
--        START_OF_PACKET_CHAR     : std_logic_vector ( 31 downto 0)  := x"060504bc"
--    );
--    port
--    (
--        -- User Interface
--        RX_DATA_IN               : in  std_logic_vector((RX_DATA_WIDTH-1) downto 0);
--        RXCTRL_IN                : in  std_logic_vector((RXCTRL_WIDTH-1) downto 0); 
--    RXENMCOMMADET_OUT        : out std_logic;
--    RXENPCOMMADET_OUT        : out std_logic;
--    RX_ENCHAN_SYNC_OUT       : out std_logic;
--    RX_CHANBOND_SEQ_IN       : in  std_logic;
--
--        -- Control Interface
--    INC_IN                   : in  std_logic; 
--    INC_OUT                  : out std_logic; 
--    PATTERN_MATCHB_OUT       : out std_logic;
--    RESET_ON_ERROR_IN        : in  std_logic;
--
--
--        -- Error Monitoring
--    ERROR_COUNT_OUT          : out std_logic_vector(7 downto 0);
--
--        -- Track Data
--    TRACK_DATA_OUT           : out std_logic;
--
--    RX_SLIDE                 : out std_logic;
--
--     
--
--        -- System Interface
--    USER_CLK                 : in std_logic;       
--    SYSTEM_RESET             : in std_logic
--);
--    end component;
--
--    component vio_0 
--        port (
--            clk : in std_logic;
--            probe_in0 : in std_logic_vector(0 downto 0);
--            probe_out0 : out std_logic_vector(0 downto 0)
--        );
--    end component;
--
--    component ila_0 
--        port (
--            clk : in std_logic;
--            probe0 : in std_logic_vector(79 downto 0);
--            probe1: in std_logic_vector(7 downto 0);
--            probe2: in std_logic_vector(0 downto 0);
--            probe3: in std_logic_vector(1 downto 0);
--            probe4: in std_logic_vector(7 downto 0);
--            probe5: in std_logic_vector(0 downto 0);
--            probe6: in std_logic_vector(0 downto 0)
--        ); 
--    end component;
--
--    component ila_1 
--        port (
--            clk : in std_logic;
--            probe0: in std_logic_vector(0 downto 0);
--            probe1: in std_logic_vector(0 downto 0)
--        ); 
--    end component;
--
----***********************************Parameter Declarations********************

  constant DLY : time := 1 ns;

--************************** Register Declarations ****************************
  attribute ASYNC_REG                          : string;
  signal gt_txfsmresetdone_r                   : std_logic;
  signal gt_txfsmresetdone_r2                  : std_logic;
  attribute ASYNC_REG of gt_txfsmresetdone_r   : signal is "TRUE";
  attribute ASYNC_REG of gt_txfsmresetdone_r2  : signal is "TRUE";
  signal gt0_txfsmresetdone_i                  : std_logic;
  signal gt0_rxfsmresetdone_i                  : std_logic;
  signal gt0_txfsmresetdone_r                  : std_logic;
  signal gt0_txfsmresetdone_r2                 : std_logic;
  attribute ASYNC_REG of gt0_txfsmresetdone_r  : signal is "TRUE";
  attribute ASYNC_REG of gt0_txfsmresetdone_r2 : signal is "TRUE";
  signal gt0_rxfsmresetdone_r                  : std_logic;
  signal gt0_rxfsmresetdone_r2                 : std_logic;
  attribute ASYNC_REG of gt0_rxfsmresetdone_r  : signal is "TRUE";
  attribute ASYNC_REG of gt0_rxfsmresetdone_r2 : signal is "TRUE";
  signal gt0_rxresetdone_r                     : std_logic;
  signal gt0_rxresetdone_r2                    : std_logic;
  signal gt0_rxresetdone_r3                    : std_logic;
  attribute ASYNC_REG of gt0_rxresetdone_r     : signal is "TRUE";
  attribute ASYNC_REG of gt0_rxresetdone_r2    : signal is "TRUE";
  attribute ASYNC_REG of gt0_rxresetdone_r3    : signal is "TRUE";



--**************************** Wire Declarations ******************************
  -------------------------- GT Wrapper Wires ------------------------------
  --________________________________________________________________________
  --________________________________________________________________________
  --GT0  (X0Y3)

  ---------------------------- Channel - DRP Ports  --------------------------
  signal gt0_drpaddr_i           : std_logic_vector(8 downto 0);
  signal gt0_drpdi_i             : std_logic_vector(15 downto 0);
  signal gt0_drpdo_i             : std_logic_vector(15 downto 0);
  signal gt0_drpen_i             : std_logic;
  signal gt0_drprdy_i            : std_logic;
  signal gt0_drpwe_i             : std_logic;
  --------------------- RX Initialization and Reset Ports --------------------
  -------------------------- RX Margin Analysis Ports ------------------------
  signal gt0_eyescandataerror_i  : std_logic;
  ------------------ Receive Ports - FPGA RX Interface Ports -----------------
  signal gt0_rxdata_i            : std_logic_vector(31 downto 0);
  ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
  signal gt0_rxcharisk_i         : std_logic_vector(3 downto 0);
  signal gt0_rxdisperr_i         : std_logic_vector(3 downto 0);
  signal gt0_rxnotintable_i      : std_logic_vector(3 downto 0);
  ------------------------ Receive Ports - RX AFE Ports ----------------------
  -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
  --signal gt0_rxslide_i           : std_logic := '0'; -- RXSLIDE_MODE = "OFF"
                                                     -- under the hood, and slide driven to 0 under the hood
  signal gt0_rxbyteisaligned_out : std_logic;
  signal gt0_rxbyterealign_out   : std_logic;
  signal gt0_rxcommadet_out      : std_logic;
  ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
  signal gt0_dmonitorout_i       : std_logic_vector(14 downto 0);
  -------------------- Receive Ports - RX Equailizer Ports -------------------
  --------------- Receive Ports - RX Fabric Output Control Ports -------------
  signal gt0_rxoutclkfabric_i    : std_logic;
  ------------- Receive Ports - RX Initialization and Reset Ports ------------
  signal gt0_rxlpmreset_i        : std_logic;
  -------------- Receive Ports -RX Initialization and Reset Ports ------------
  signal gt0_rxresetdone_i       : std_logic;
  --------------------- TX Initialization and Reset Ports --------------------
  ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
  signal gt0_txdata_i            : std_logic_vector(31 downto 0);
  ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
  signal gt0_txcharisk_i         : std_logic_vector(3 downto 0);
  --------------- Transmit Ports - TX Configurable Driver Ports --------------
  ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
  signal gt0_txoutclkfabric_i    : std_logic;
  signal gt0_txoutclkpcs_i       : std_logic;
  ------------- Transmit Ports - TX Initialization and Reset Ports -----------
  signal gt0_txresetdone_i       : std_logic;



  --____________________________COMMON PORTS________________________________
  -------------------------- Common Block - PLL Ports ------------------------
  signal gt0_pll0lock_i       : std_logic;
  signal gt0_pll0refclklost_i : std_logic;
  signal gt0_pll0reset_i      : std_logic;



  ------------------------------- Global Signals -----------------------------
  signal gt0_tx_system_reset_c : std_logic;
  signal gt0_rx_system_reset_c : std_logic;
  signal tied_to_ground_i      : std_logic;
  signal tied_to_ground_vec_i  : std_logic_vector(63 downto 0);
  signal tied_to_vcc_i         : std_logic;
  signal tied_to_vcc_vec_i     : std_logic_vector(7 downto 0);



  attribute keep         : string;
  ------------------------------- User Clocks ---------------------------------
  signal gt0_txusrclk_i  : std_logic;
  signal gt0_txusrclk2_i : std_logic;
  signal gt0_rxusrclk_i  : std_logic;
  signal gt0_rxusrclk2_i : std_logic;

  signal gt0_txmmcm_lock_i  : std_logic;
  signal gt0_rxmmcm_lock_i  : std_logic;


  ----------------------------- Reference Clocks ----------------------------


  ----------------------- Frame check/gen Module Signals --------------------

  signal gt0_matchn_i            : std_logic;
  signal gt0_track_data_i        : std_logic;
  signal gt0_error_count_i       : std_logic_vector(7 downto 0);
  signal gt0_frame_check_reset_i : std_logic;
  signal gt0_inc_in_i            : std_logic;
  signal gt0_inc_out_i           : std_logic;

  signal reset_on_data_error_i : std_logic;
  signal track_data_out_i      : std_logic;
  signal track_data_out_ila_i  : std_logic_vector(0 downto 0);

  ----------------------- Chipscope Signals ---------------------------------



  signal zero_vector_rx_80    : std_logic_vector ((80 -32) -1 downto 0) := (others => '0');
  signal zero_vector_rx_8     : std_logic_vector ((8 -4) -1 downto 0)   := (others => '0');
  signal gt0_rxdata_ila       : std_logic_vector (79 downto 0);
  signal gt0_rxdatavalid_ila  : std_logic_vector (1 downto 0);
  signal gt0_rxcharisk_ila    : std_logic_vector (7 downto 0);
  signal gt0_txmmcm_lock_ila  : std_logic_vector (0 downto 0);
  signal gt0_rxmmcm_lock_ila  : std_logic_vector (0 downto 0);
  signal gt0_rxresetdone_ila  : std_logic_vector (0 downto 0);
  signal gt0_txresetdone_ila  : std_logic_vector (0 downto 0);
  signal tied_to_ground_ila_i : std_logic_vector (0 downto 0);
  -- update with the actual reset name
  signal soft_reset_i         : std_logic;
  signal soft_reset_vio_i     : std_logic_vector (0 downto 0);
  signal gt0_rxfsmresetdone_s : std_logic_vector(0 downto 0);


  function and_reduce(arg : std_logic_vector) return std_logic is
    variable result : std_logic;
  begin
    result := '1';
    for i in arg'range loop
      result := result and arg(i);
    end loop;
    return result;
  end;

  signal probe0_unpack_telemetry : std_logic_vector(7 downto 0);
  signal probe0 : std_logic_vector(7 downto 0);
  signal probe1 : std_logic_vector(7 downto 0);
  signal probe2 : std_logic_vector(7 downto 0);
  signal probe3 : std_logic_vector(7 downto 0);
  signal probe4 : std_logic_vector(7 downto 0);
  signal probe5 : std_logic_vector(7 downto 0);
  signal probe6 : std_logic_vector(7 downto 0);
  signal probe7 : std_logic_vector(7 downto 0);

  signal probe0_rx : std_logic_vector(7 downto 0);
  signal probe1_rx : std_logic_vector(7 downto 0);
  signal probe2_rx : std_logic_vector(7 downto 0);
  signal probe3_rx : std_logic_vector(7 downto 0);
  signal probe4_rx : std_logic_vector(7 downto 0);
  signal probe5_rx : std_logic_vector(7 downto 0);
  signal probe6_rx : std_logic_vector(7 downto 0);
  signal probe7_rx : std_logic_vector(7 downto 0);

-- telemetry

  signal clk_128M   : std_logic;
  signal soft_reset_cnt : std_logic_vector(15 downto 0) := (others=>'0');
  signal soft_reset_auto : std_logic := '0';

--  signal vio_slide           : std_logic;
--  signal vio_slide_ila           : std_logic_vector(0 downto 0);

--  signal r_vio_slide : std_logic := '0';
--  signal r_vio_slide_pulse : std_logic := '0';
--  signal gt0_rxslide_i2 : std_logic := '0';

--**************************** Main Body of Code *******************************
begin

  --  Static signal Assigments
  tied_to_ground_i     <= '0';
  tied_to_ground_vec_i <= x"0000000000000000";
  tied_to_vcc_i        <= '1';
  tied_to_vcc_vec_i    <= "11111111";

  
  -- outputs
  data_out <= gt0_rxdata_i;
  DATA_CLK_OUT <= gt0_rxusrclk2_i;
  data_is_k_out <= gt0_rxcharisk_i;
  SOFT_RESET_OUT <= soft_reset_i;
  ----------------------------- The GT Wrapper -----------------------------

  -- Use the instantiation template in the example directory to add the GT wrapper to your design.
  -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
  -- checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
  -- enabled, bonding should occur after alignment
  -- While connecting the GT TX/RX Reset ports below, please add a delay of
  -- minimum 500ns as mentioned in AR 43482.

  -- was in: rtl/gt_ip/gt_serial_telem_rx.vhd, now generated by xci and not committed to version control
  gt_serial_telem_rx_i : entity work.gt_serial_telem_rx
    port map
    (
      soft_reset_tx_in            => soft_reset_i,
      soft_reset_rx_in            => soft_reset_i,
      DONT_RESET_ON_DATA_ERROR_IN => tied_to_vcc_i,
      Q0_CLK1_GTREFCLK_PAD_N_IN   => Q0_CLK1_GTREFCLK_PAD_N_IN,
      Q0_CLK1_GTREFCLK_PAD_P_IN   => Q0_CLK1_GTREFCLK_PAD_P_IN,
      GT0_TX_MMCM_LOCK_OUT        => gt0_txmmcm_lock_i,
      GT0_RX_MMCM_LOCK_OUT        => gt0_rxmmcm_lock_i,
      GT0_TX_FSM_RESET_DONE_OUT   => gt0_txfsmresetdone_i,
      GT0_RX_FSM_RESET_DONE_OUT   => gt0_rxfsmresetdone_i,
      GT0_DATA_VALID_IN           => gt0_track_data_i,

      GT0_TXUSRCLK_OUT  => gt0_txusrclk_i,
      GT0_TXUSRCLK2_OUT => gt0_txusrclk2_i,
      GT0_RXUSRCLK_OUT  => gt0_rxusrclk_i,
      GT0_RXUSRCLK2_OUT => gt0_rxusrclk2_i,

      --_____________________________________________________________________
      --_____________________________________________________________________
      --GT0  (X0Y3)

      ---------------------------- Channel - DRP Ports  --------------------------
      gt0_drpaddr_in           => gt0_drpaddr_i,
      gt0_drpdi_in             => gt0_drpdi_i,
      gt0_drpdo_out            => gt0_drpdo_i,
      gt0_drpen_in             => gt0_drpen_i,
      gt0_drprdy_out           => gt0_drprdy_i,
      gt0_drpwe_in             => gt0_drpwe_i,
      --------------------- RX Initialization and Reset Ports --------------------
      gt0_eyescanreset_in      => tied_to_ground_i,
      gt0_rxuserrdy_in         => tied_to_vcc_i,
      -------------------------- RX Margin Analysis Ports ------------------------
      gt0_eyescandataerror_out => gt0_eyescandataerror_i,
      gt0_eyescantrigger_in    => tied_to_ground_i,
      ------------------ Receive Ports - FPGA RX Interface Ports -----------------
      gt0_rxdata_out           => gt0_rxdata_i,
      ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
      gt0_rxcharisk_out        => gt0_rxcharisk_i,
      gt0_rxdisperr_out        => gt0_rxdisperr_i,
      gt0_rxnotintable_out     => gt0_rxnotintable_i,
      ------------------------ Receive Ports - RX AFE Ports ----------------------
      gt0_gtprxn_in            => RXN_IN,
      gt0_gtprxp_in            => RXP_IN,
      -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
      gt0_rxbyteisaligned_out  => gt0_rxbyteisaligned_out,
      gt0_rxbyterealign_out    => gt0_rxbyterealign_out,
      gt0_rxcommadet_out       => gt0_rxcommadet_out,
      --gt0_rxslide_in           => gt0_rxslide_i,
--# https://support.xilinx.com/s/article/67147?language=en_US
--You should uncheck RXSLIDE and manually check RXPCOMMAALIGNEN and RXMCOMMAALIGNEN if comma alignment is to be used.
--If this is not done, RXPCOMMAALIGNEN and RXMCOMMAALIGNEN will be tied to ground and comma alignment will not work.

      gt0_rxmcommaalignen_in   => '1',
      gt0_rxpcommaalignen_in   => '1',

      ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
      gt0_dmonitorout_out      => gt0_dmonitorout_i,
      -------------------- Receive Ports - RX Equailizer Ports -------------------
      gt0_rxlpmhfhold_in       => tied_to_ground_i,
      gt0_rxlpmlfhold_in       => tied_to_ground_i,
      --------------- Receive Ports - RX Fabric Output Control Ports -------------
      gt0_rxoutclkfabric_out   => gt0_rxoutclkfabric_i,
      ------------- Receive Ports - RX Initialization and Reset Ports ------------
      gt0_gtrxreset_in         => tied_to_ground_i,
      gt0_rxlpmreset_in        => gt0_rxlpmreset_i,
      -------------- Receive Ports -RX Initialization and Reset Ports ------------
      gt0_rxresetdone_out      => gt0_rxresetdone_i,
      --------------------- TX Initialization and Reset Ports --------------------
      gt0_gttxreset_in         => tied_to_ground_i,
      gt0_txuserrdy_in         => tied_to_vcc_i,
      ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
      gt0_txdata_in            => gt0_txdata_i,
      ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
      gt0_txcharisk_in         => gt0_txcharisk_i,
      --------------- Transmit Ports - TX Configurable Driver Ports --------------
      gt0_gtptxn_out           => TXN_OUT,
      gt0_gtptxp_out           => TXP_OUT,
      ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
      gt0_txoutclkfabric_out   => gt0_txoutclkfabric_i,
      gt0_txoutclkpcs_out      => gt0_txoutclkpcs_i,
      ------------- Transmit Ports - TX Initialization and Reset Ports -----------
      gt0_txresetdone_out      => gt0_txresetdone_i,



      --____________________________COMMON PORTS________________________________
      GT0_PLL0RESET_OUT      => open,
      GT0_PLL0OUTCLK_OUT     => open,
      GT0_PLL0OUTREFCLK_OUT  => open,
      GT0_PLL0LOCK_OUT       => open,
      GT0_PLL0REFCLKLOST_OUT => open,
      GT0_PLL1OUTCLK_OUT     => open,
      GT0_PLL1OUTREFCLK_OUT  => open,
      gt0_rxpolarity_in      => '0',
      sysclk_in              => clk_128M -- DRP_CLK_IN
      );

  -- IBUFDS_DRP_CLK : IBUFDS
  -- port map
  --   (
  --      I  => DRP_CLK_IN_P,
  --      IB => DRP_CLK_IN_N,
  --      O  => DRPCLK_IN
  --   );

  -- DRP_CLK_BUFG : BUFG 
  -- port map 
  --  (
  --      I    => DRPCLK_IN,
  --      O    => drpclk_in_i 
  --  );

  clk_128M <= DRP_CLK_IN;


  -------------------------- User Module Resets -----------------------------
  -- All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
  -- are held in reset till the RESETDONE goes high. 
  -- The RESETDONE is registered a couple of times on USRCLK2 and connected 
  -- to the reset of the modules

  process(gt0_rxusrclk2_i, gt0_rxresetdone_i)
  begin
    if(gt0_rxresetdone_i = '0') then
      gt0_rxresetdone_r  <= '0' after DLY;
      gt0_rxresetdone_r2 <= '0' after DLY;
      gt0_rxresetdone_r3 <= '0' after DLY;
    elsif (gt0_rxusrclk2_i'event and gt0_rxusrclk2_i = '1') then
      gt0_rxresetdone_r  <= gt0_rxresetdone_i  after DLY;
      gt0_rxresetdone_r2 <= gt0_rxresetdone_r  after DLY;
      gt0_rxresetdone_r3 <= gt0_rxresetdone_r2 after DLY;
    end if;
  end process;

  process(gt0_txusrclk2_i, gt0_txfsmresetdone_i)
  begin
    if(gt0_txfsmresetdone_i = '0') then
      gt0_txfsmresetdone_r  <= '0' after DLY;
      gt0_txfsmresetdone_r2 <= '0' after DLY;
    elsif (gt0_txusrclk2_i'event and gt0_txusrclk2_i = '1') then
      gt0_txfsmresetdone_r  <= gt0_txfsmresetdone_i after DLY;
      gt0_txfsmresetdone_r2 <= gt0_txfsmresetdone_r after DLY;
    end if;
  end process;


  ------------------------------ Frame Generators ---------------------------
  -- The example design uses Block RAM based frame generators to provide test
  -- data to the GTs for transmission. By default the frame generators are 
  -- loaded with an incrementing data sequence that includes commas/alignment
  -- characters for alignment. If your protocol uses channel bonding, the 
  -- frame generator will also be preloaded with a channel bonding sequence.

  -- You can modify the data transmitted by changing the INIT values of the frame
  -- generator in this file. Pay careful attention to bit order and the spacing
  -- of your control and alignment characters.

--  gt0_frame_gen : entity work.gt_serial_telem_rx_GT_FRAME_GEN
--    generic map
--    (
--      WORDS_IN_BRAM => EXAMPLE_WORDS_IN_BRAM
--      )
--    port map
--    (
--      -- User Interface
--      TX_DATA_OUT(79 downto 48) => gt0_txdata_float_i,
--      TX_DATA_OUT(15 downto 0)  => gt0_txdata_float16_i,
--      TX_DATA_OUT(47 downto 16) => gt0_txdata_i,
-- 
--      TXCTRL_OUT(7 downto 4) => gt0_txcharisk_float_i,
--      TXCTRL_OUT(3 downto 0) => gt0_txcharisk_i,
--      -- System Interface
--      USER_CLK               => gt0_txusrclk2_i,
--      SYSTEM_RESET           => gt0_tx_system_reset_c
--      );

  ---------------------------------- Frame Checkers -------------------------
  -- The example design uses Block RAM based frame checkers to verify incoming  
  -- data. By default the frame generators are loaded with a data sequence that 
  -- matches the outgoing sequence of the frame generators for the TX ports.

  -- You can modify the expected data sequence by changing the INIT values of the frame
  -- checkers in this file. Pay careful attention to bit order and the spacing
  -- of your control and alignment characters.

  -- When the frame checker receives data, it attempts to synchronise to the 
  -- incoming pattern by looking for the first sequence in the pattern. Once it 
  -- finds the first sequence, it increments through the sequence, and indicates an 
  -- error whenever the next value received does not match the expected value.

  gt0_frame_check_reset_i <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES = 0) else gt0_matchn_i;

  -- gt0_frame_check0 is always connected to the lane with the start of char 
  -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
  gt0_inc_in_i <= '0';

--  gt0_frame_check : entity work.gt_serial_telem_rx_GT_FRAME_CHECK
--    generic map
--    (
--      RX_DATA_WIDTH        => 32,
--      RXCTRL_WIDTH         => 4,
--      COMMA_DOUBLE         => x"bcbc",
--      WORDS_IN_BRAM        => EXAMPLE_WORDS_IN_BRAM,
--      START_OF_PACKET_CHAR => x"bcbcbcbc"
--      )
--    port map
--    (
--      -- GT Interface
--      RX_DATA_IN         => gt0_rxdata_i,
--      RXCTRL_IN          => gt0_rxcharisk_i,
--      RXENMCOMMADET_OUT  => open,
--      RXENPCOMMADET_OUT  => open,
--      RX_ENCHAN_SYNC_OUT => open,
--      RX_CHANBOND_SEQ_IN => tied_to_ground_i,
--      -- Control Interface
--      INC_IN             => gt0_inc_in_i,
--      INC_OUT            => gt0_inc_out_i,
--      PATTERN_MATCHB_OUT => gt0_matchn_i,
--      RESET_ON_ERROR_IN  => gt0_frame_check_reset_i,
--      -- System Interface
--      USER_CLK           => gt0_rxusrclk2_i,
--      SYSTEM_RESET       => gt0_rx_system_reset_c,
--      ERROR_COUNT_OUT    => gt0_error_count_i,
--      RX_SLIDE           => gt0_rxslide_i,
--      TRACK_DATA_OUT     => gt0_track_data_i
--      );




--  TRACK_DATA_OUT <= track_data_out_i;

  track_data_out_i <=
    gt0_track_data_i;



--  probe0_unpack_telemetry <= "00" & r_sticky_led_out & okay_led_out & r_sticky_pll2_locked & r_sticky_pll_locked & '0' & pll_locked;
--  gen_debug : if g_debug = '1' generate
--
--    inst_ila_8x8_0 : entity work.ila_8x8
--      port map (
--        clk    => clk_256M,
--        probe0 => probe0_unpack_telemetry,
--        probe1 => "00000000",
--        probe2 => "00000000",
--        probe3 => "00000000",
--        probe4 => "00000000",
--        probe5 => "00000000",
--        probe6 => "00000000",
--        probe7 => "00000000"
--        );
--  end generate gen_debug;



-------------------------------------------------------------------------------
----------------------------- Debug Signals assignment -----------------------

------------ optional Ports assignments --------------
------------------------------------------------------ 

  -- assign resets for frame_gen modules
  gt0_tx_system_reset_c <= not gt0_txfsmresetdone_r2;

  -- assign resets for frame_check modules
  gt0_rx_system_reset_c <= not gt0_rxresetdone_r3;


  gt0_rxlpmreset_i <= '0';
  gt0_drpaddr_i    <= (others => '0');
  gt0_drpdi_i      <= (others => '0');
  gt0_drpen_i      <= '0';
  gt0_drpwe_i      <= '0';


  tied_to_ground_ila_i(0) <= '0';
  gt0_rxfsmresetdone_s(0) <= gt0_rxfsmresetdone_i;

  soft_reset_i <= soft_reset_auto or soft_reset_vio_i(0);

  no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate
      soft_reset_vio_i <= (others=>'0');
  end generate no_chipscope;

  chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate
    -- vio core insertion for driving soft_reset_i
      vio_gt_inst : entity work.vio_0 port map (
        clk        => clk_128M,  -- input DRP_CLK_IN
        probe_in0  => gt0_rxfsmresetdone_s,
        probe_out0 => soft_reset_vio_i
        );
  end generate chipscope;


  process(clk_128M)begin
      if rising_edge(clk_128M) then
          if(rst_128M='1')then
              soft_reset_auto <= '1';
              soft_reset_cnt <= (others=>'0');
          elsif(soft_reset_cnt=X"FFFF")then
              soft_reset_auto <= '0';
          else
              soft_reset_cnt <= soft_reset_cnt + '1';
          end if;
      end if;
  end process;

  -- xilinx doesn't need this, but modelim errors out with:
  -- Signal "vio_slide" is type ieee.std_logic_1164.STD_LOGIC; expecting type ieee.std_logic_1164.STD_LOGIC_VECTOR.
--  vio_slide_ila(0) <= vio_slide; 

--  vio_gt_slip_inst : entity work.vio_0 port map (
--    clk        => gt0_rxusrclk2_i,  -- input clk
--    probe_in0  => gt0_rxfsmresetdone_s,
--    probe_out0 => vio_slide_ila
--    );

--  proc_cnt_input : process(gt0_rxusrclk2_i)
--  begin
--    if rising_edge(gt0_rxusrclk2_i) then
--      r_vio_slide <= vio_slide;
--      r_vio_slide_pulse <= vio_slide and not r_vio_slide; -- rising edge detect
--      gt0_rxslide_i2 <= gt0_rxslide_i or r_vio_slide_pulse;      
--    end if;
--  end process;


  gt0_rxdata_ila <= zero_vector_rx_80 & gt0_rxdata_i;

  gt0_rxdatavalid_ila(0) <= '0';
  gt0_rxdatavalid_ila(1) <= '0';

  gt0_rxcharisk_ila <= zero_vector_rx_8 & gt0_rxcharisk_i;


  gt0_txmmcm_lock_ila(0) <= gt0_txmmcm_lock_i;

  gt0_rxmmcm_lock_ila(0) <= gt0_rxmmcm_lock_i;
  gt0_rxresetdone_ila(0) <= gt0_rxresetdone_i;
  gt0_txresetdone_ila(0) <= gt0_txresetdone_i;

  track_data_out_ila_i(0) <= track_data_out_i;


-- ila core insertion for observing data and control signals
  ila_tx0_inst : entity work.ila_1 port map (
    clk    => gt0_txusrclk_i,  -- input clk
    probe0 => gt0_txmmcm_lock_ila,
    probe1 => gt0_txresetdone_ila
    );

  ila_rx0_inst : entity work.ila_gt_rx_0 port map (
    clk    => gt0_rxusrclk_i,  -- input clk
    probe0 => gt0_rxdata_ila,
    probe1 => gt0_error_count_i,
    probe2 => track_data_out_ila_i,
    probe3 => gt0_rxdatavalid_ila,
    probe4 => gt0_rxcharisk_ila,
    probe5 => gt0_rxmmcm_lock_ila,
    probe6 => gt0_rxresetdone_ila
    );






  probe0 <= "0" & gt0_rxmmcm_lock_ila(0) & gt0_rxresetdone_ila(0) & track_data_out_ila_i(0) &
            gt0_rxresetdone_ila(0) & gt0_rxcommadet_out & gt0_rxbyterealign_out & gt0_rxbyteisaligned_out;
  probe1 <= gt0_error_count_i;
  probe2 <= gt0_rxcharisk_ila;
  probe3 <= "00000"  & gt0_frame_check_reset_i &gt0_matchn_i & gt0_inc_out_i;
  probe4 <= "00000000";
  probe5 <= "00000000";
  probe6 <= "00000000";
  probe7 <= "00000000";
  
  ila_8x8_inst : entity work.ila_8x8 port map (
    clk    => gt0_txusrclk_i,
    probe0 => probe0,
    probe1 => probe1,
    probe2 => probe2,
    probe3 => probe3,
    probe4 => probe4,
    probe5 => probe5,
    probe6 => probe6,
    probe7 => probe7
    );


  probe0_rx <= "0" & gt0_rxmmcm_lock_ila(0) & gt0_rxresetdone_ila(0) & track_data_out_ila_i(0) &
            gt0_rxresetdone_ila(0) & gt0_rxcommadet_out & gt0_rxbyterealign_out & gt0_rxbyteisaligned_out;
  probe1_rx <= gt0_error_count_i;
  probe2_rx <= gt0_rxcharisk_ila;
  probe3_rx <= "00000" & gt0_frame_check_reset_i &gt0_matchn_i & gt0_inc_out_i;
  probe4_rx <= gt0_rxnotintable_i & gt0_rxdisperr_i;
  probe5_rx <= "00000000";
  probe6_rx <= "00000000";
  probe7_rx <= "00000000";
  ila_8x8_rx_inst : entity work.ila_8x8 port map (
    clk    => gt0_rxusrclk_i,
    probe0 => probe0_rx,
    probe1 => probe1_rx,
    probe2 => probe2_rx,
    probe3 => probe3_rx,
    probe4 => probe4_rx,
    probe5 => probe5_rx,
    probe6 => probe6_rx,
    probe7 => probe7_rx 
    );

  

end RTL;


