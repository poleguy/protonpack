do not use 